package filter_pkg;
typedef struct packed {
	logic dummy;
}filter_to_pad_t;

typedef struct packed{
	logic dummy;
}pad_to_filter_t;
endpackage